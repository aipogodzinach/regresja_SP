��e,      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.1�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�P1��P2��P3��P4��P5��P6�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        h@KhAKhBh(h+K ��h-��R�(KK��h2�f8�����R�(KhJNNNJ����J����K t�b�C              �?�t�bhNh&�scalar���hIC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hI�C       �t�bK��R�}�(hK�
node_count�K�nodes�h(h+K ��h-��R�(KK��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hzh2�i8�����R�(KhJNNNJ����J����K t�bK ��h{h�K��h|h�K��h}hZK��h~hZK ��hh�K(��h�hZK0��uK8KKt�b�Bh         
                    @�8��8��?             H@       	                    @8�Z$���?             :@                           @      �?              @                           @      �?             @������������������������       �                     �?������������������������       �                     @                           @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@������������������������       �                     6@�t�b�values�h(h+K ��h-��R�(KKKK��hZ�C�      @      F@      @      6@      @      @      �?      @      �?                      @      @      �?      @                      �?              2@              6@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        h@KhAKhBh(h+K ��h-��R�(KK��hZ�C              �?�t�bhNh_hIC       ���R�hcKhdhgKh(h+K ��h-��R�(KK��hI�C       �t�bK��R�}�(hKhqK	hrh(h+K ��h-��R�(KK	��hy�B�                             @      �?!             H@                           @d}h���?             ,@������������������������       �                     �?                           @8�Z$���?             *@                           @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     A@�t�bh�h(h+K ��h-��R�(KK	KK��hZ�C�      @     �F@      @      &@      �?               @      &@       @      �?              �?       @                      $@              A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        h@KhAKhBh(h+K ��h-��R�(KK��hZ�C              �?�t�bhNh_hIC       ���R�hcKhdhgKh(h+K ��h-��R�(KK��hI�C       �t�bK��R�}�(hKhqK	hrh(h+K ��h-��R�(KK	��hy�B�                             @      �?             H@������������������������       �                     @                           @���7�?             F@                           @z�G�z�?             $@                           @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     A@�t�bh�h(h+K ��h-��R�(KK	KK��hZ�C�      @      E@      @               @      E@       @       @       @      �?              �?       @                      @              A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        h@KhAKhBh(h+K ��h-��R�(KK��hZ�C              �?�t�bhNh_hIC       ���R�hcKhdhgKh(h+K ��h-��R�(KK��hI�C       �t�bK��R�}�(hKhqKhrh(h+K ��h-��R�(KK��hy�Bh                             @�q�q��?             H@                           @����X�?             ,@                           @�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �                     @       
                     @г�wY;�?             A@       	                    @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     <@�t�bh�h(h+K ��h-��R�(KKKK��hZ�C�      &@     �B@      $@      @      $@      �?              �?      $@                      @      �?     �@@      �?      @              @      �?                      <@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        h@KhAKhBh(h+K ��h-��R�(KK��hZ�C              �?�t�bhNh_hIC       ���R�hcKhdhgKh(h+K ��h-��R�(KK��hI�C       �t�bK��R�}�(hKhqKhrh(h+K ��h-��R�(KK��hy�Bh                              @�8��8��?#             H@                           @      �?	             (@������������������������       �                      @                           @ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?       
                    @������?             B@       	                    @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     ?@�t�bh�h(h+K ��h-��R�(KKKK��hZ�C�      @      F@      @      "@       @              �?      "@              "@      �?              �?     �A@      �?      @      �?                      @              ?@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        h@KhAKhBh(h+K ��h-��R�(KK��hZ�C              �?�t�bhNh_hIC       ���R�hcKhdhgKh(h+K ��h-��R�(KK��hI�C       �t�bK��R�}�(hKhqKhrh(h+K ��h-��R�(KK��hy�Bh                             @ �q�q�?             H@                           @�q�q�?             @������������������������       �                     �?                            @      �?              @������������������������       �                     �?������������������������       �                     �?       
                    @����?�?            �F@       	                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �E@�t�bh�h(h+K ��h-��R�(KKKK��hZ�C�       @      G@      �?       @              �?      �?      �?              �?      �?              �?      F@      �?      �?              �?      �?                     �E@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        h@KhAKhBh(h+K ��h-��R�(KK��hZ�C              �?�t�bhNh_hIC       ���R�hcKhdhgKh(h+K ��h-��R�(KK��hI�C       �t�bK��R�}�(hK hqKhrh(h+K ��h-��R�(KK��hy�C8������������������������       �                     H@�t�bh�h(h+K ��h-��R�(KKKK��hZ�C              H@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        h@KhAKhBh(h+K ��h-��R�(KK��hZ�C              �?�t�bhNh_hIC       ���R�hcKhdhgKh(h+K ��h-��R�(KK��hI�C       �t�bK��R�}�(hKhqKhrh(h+K ��h-��R�(KK��hy�B�                             @r�q��?             H@������������������������       �                     @                           @�C��2(�?             F@                           @�<ݚ�?             "@������������������������       �                     @                           @�q�q�?             @������������������������       �                      @������������������������       �                     �?	                           @ >�֕�?            �A@
                           @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     >@�t�bh�h(h+K ��h-��R�(KKKK��hZ�C�       @      D@      @              @      D@       @      @              @       @      �?       @                      �?       @     �@@       @      @              @       @                      >@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        h@KhAKhBh(h+K ��h-��R�(KK��hZ�C              �?�t�bhNh_hIC       ���R�hcKhdhgKh(h+K ��h-��R�(KK��hI�C       �t�bK��R�}�(hKhqKhrh(h+K ��h-��R�(KK��hy�Bh                             @8��8���?             H@                           @      �?             @                           @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @       
                    @���N8�?             E@       	                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �C@�t�bh�h(h+K ��h-��R�(KKKK��hZ�C�      @     �E@      @      @      @      �?      @                      �?               @       @      D@       @      �?              �?       @                     �C@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        h@KhAKhBh(h+K ��h-��R�(KK��hZ�C              �?�t�bhNh_hIC       ���R�hcKhdhgKh(h+K ��h-��R�(KK��hI�C       �t�bK��R�}�(hKhqKhrh(h+K ��h-��R�(KK��hy�Bh                             @      �?             H@                           @�q�q�?             @������������������������       �                      @������������������������       �                     �?       
                    @����?�?            �F@                           @r�q��?             @������������������������       �                      @       	                    @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                    �C@�t�bh�h(h+K ��h-��R�(KKKK��hZ�C�      @     �F@       @      �?       @                      �?      �?      F@      �?      @               @      �?      @      �?                      @             �C@�t�bubhhubehhub.